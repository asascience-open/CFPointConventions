netcdf trajectoryProfile-Multidimensional-MultipleTrajectories-H.6.1 {
dimensions:
	trajectory = UNLIMITED ; // (6 currently)
	profile = 10 ;
	z = 8 ;
variables:
	float lat(trajectory, profile) ;
		lat:units = "degrees_north" ;
		lat:long_name = "Latitude" ;
		lat:standard_name = "latitude" ;
		lat:missing_value = -999.9f ;
	float lon(trajectory, profile) ;
		lon:units = "degrees_east" ;
		lon:long_name = "Longitude" ;
		lon:standard_name = "longitude" ;
		lon:missing_value = -999.9f ;
	int trajectory(trajectory) ;
		trajectory:cf_role = "trajectory_id" ;
	float alt(trajectory, profile, z) ;
		alt:standard_name = "altitude" ;
		alt:long_name = "height below mean sea level" ;
		alt:units = "m" ;
		alt:positive = "down" ;
		alt:axis = "Z" ;
		alt:missing_value = -999.f ;
	int time(trajectory, profile) ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
		time:missing_value = -999 ;
	float temperature(trajectory, profile, z) ;
		temperature:long_name = "Water Temperature" ;
		temperature:standard_name = "air_temperature" ;
		temperature:units = "Celsius" ;
		temperature:coordinates = "time lat lon alt" ;
		temperature:missing_value = -999.9f ;
	float salinity(trajectory, profile, z) ;
		salinity:long_name = "Sea Water Salinity" ;
		salinity:standard_name = "sea_water_salinity" ;
		salinity:units = "PSU" ;
		salinity:coordinates = "time lat lon alt" ;
		salinity:missing_value = -999.9f ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:featureType = "trajectoryProfile" ;
}
