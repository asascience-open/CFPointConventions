netcdf profile-Incomplete-MultiDimensional-MultipleProfiles-H.3.2 {
dimensions:
	profile = 142 ;
	alt = 42 ;
variables:
	float lat(profile) ;
		lat:units = "degrees_north" ;
		lat:long_name = "station latitude" ;
		lat:standard_name = "latitude" ;
	float lon(profile) ;
		lon:units = "degrees_east" ;
		lon:long_name = "station longitude" ;
		lon:standard_name = "longitude" ;
	int profile(profile) ;
		profile:cf_role = "profile_id" ;
	int time(profile) ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
	float alt(profile, alt) ;
		alt:units = "m" ;
		alt:standard_name = "altitude" ;
		alt:long_name = "height above mean sea level" ;
		alt:positive = "up" ;
		alt:axis = "Z" ;
	float temperature(profile, alt) ;
		temperature:long_name = "Air Temperature" ;
		temperature:units = "Celsius" ;
		temperature:coordinates = "time lat lon alt" ;
	float humidity(profile, alt) ;
		humidity:long_name = "Humidity" ;
		humidity:standard_name = "specific_humidity" ;
		humidity:units = "Percent" ;
		humidity:coordinates = "time lat lon alt" ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:featureType = "profile" ;
}
