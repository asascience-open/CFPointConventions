netcdf timeSeriesProfile-Ragged-SingeStation-9.5.3 {
dimensions:
	profile = 4 ;
	obs = 10 ;
	name_strlen = 50 ;
variables:
	double lat ;
		lat:units = "degrees_north" ;
		lat:long_name = "station latitude" ;
		lat:standard_name = "latitude" ;
	double lon ;
		lon:units = "degrees_east" ;
		lon:long_name = "station longitude" ;
		lon:standard_name = "longitude" ;
	int station_info ;
		station_info:long_name = "station info" ;
	char station_name(name_strlen) ;
		station_name:cf_role = "timeseries_id" ;
		station_name:long_name = "station name" ;
	int profile(profile) ;
		profile:cf_role = "profile_id" ;
	int time(profile) ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
	int row_size(profile) ;
		row_size:long_name = "number of obs in this profile" ;
		row_size:sample_dimension = "obs" ;
	double height(obs) ;
		height:long_name = "height above sea surface" ;
		height:standard_name = "height" ;
		height:units = "meters" ;
		height:axis = "Z" ;
		height:positive = "up" ;
	double temperature(obs) ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:long_name = "Water Temperature" ;
		temperature:units = "Celsius" ;
		temperature:coordinates = "time lat lon height" ;

// global attributes:
		:CF\:featureType = "timeSeriesProfile" ;
}
