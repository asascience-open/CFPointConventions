netcdf timeSeries-Incomplete-MultiDimensional-MultipleStations-H.2.2 {
dimensions:
	station = UNLIMITED ; // (10 currently)
	obs = 20 ;
	name_strlen = 50 ;
variables:
	float lat(station) ;
		lat:units = "degrees_north" ;
		lat:long_name = "station latitude" ;
		lat:standard_name = "latitude" ;
	float lon(station) ;
		lon:units = "degrees_east" ;
		lon:long_name = "station longitude" ;
		lon:standard_name = "longitude" ;
	float station_elevation(station) ;
		station_elevation:long_name = "height above the geoid" ;
		station_elevation:standard_name = "surface_altitude" ;
		station_elevation:units = "m" ;
	int station_info(station) ;
		station_info:long_name = "station info" ;
	char station_name(station, name_strlen) ;
		station_name:cf_role = "timeseries_id" ;
		station_name:long_name = "station name" ;
	float alt(station) ;
		alt:long_name = "vertical distance above the surface" ;
		alt:standard_name = "height" ;
		alt:units = "m" ;
		alt:positive = "up" ;
		alt:axis = "Z" ;
	int time(station, obs) ;
		time:long_name = "time of measurement" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
		time:missing_value = -999 ;
	float temperature(station, obs) ;
		temperature:long_name = "Air Temperature" ;
		temperature:standard_name = "air_temperature" ;
		temperature:units = "Celsius" ;
		temperature:coordinates = "time lat lon alt" ;
		temperature:missing_value = -999.9f ;
	float humidity(station, obs) ;
		humidity:long_name = "Humidity" ;
		humidity:standard_name = "specific_humidity" ;
		humidity:units = "Percent" ;
		humidity:coordinates = "time lat lon alt" ;
		humidity:missing_value = -999.9f ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:featureType = "timeSeries" ;
}
