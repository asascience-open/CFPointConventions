netcdf profile-Orthogonal-SingleDimensional-SingleProfile-H.3.3 {
dimensions:
	z = 42 ;
variables:
	float lat ;
		lat:units = "degrees_north" ;
		lat:long_name = "station latitude" ;
		lat:standard_name = "latitude" ;
	float lon ;
		lon:units = "degrees_east" ;
		lon:long_name = "station longitude" ;
		lon:standard_name = "longitude" ;
	int profile ;
		profile:cf_role = "profile_id" ;
	int time ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
	float z(z) ;
		z:units = "m" ;
		z:standard_name = "altitude" ;
		z:long_name = "height above mean sea level" ;
		z:positive = "up" ;
		z:axis = "Z" ;
	float temperature(z) ;
		temperature:long_name = "Water Temperature" ;
		temperature:units = "Celsius" ;
		temperature:coordinates = "time lat lon z" ;
	float humidity(z) ;
		humidity:long_name = "Humidity" ;
		humidity:standard_name = "specific_humidity" ;
		humidity:units = "Percent" ;
		humidity:coordinates = "time lat lon z" ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:featureType = "profile" ;
}
